module master (
    input          i_clk,
    input          i_rstn,
    output         o_valid,
    input          i_ready,
    output  [31:0] o_data,
    input   [31:0] i_data
);

endmodule

