module top (
	input				i_CLK_top,
	input				i_RESETn_top,
	input	[31:0]		i_i_DATA_top,
	output	[31:0]		o_o_DATA_top,
);
endmoduleHello