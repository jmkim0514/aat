module top (
	input				i_CLK_top,
	input				i_RESETn_top,
	input	[31:0]		i_DATA_top,
	output	[31:0]		o_DATA_top,
);
endmodule