
module slave (
    input          i_clk,
    input          i_rstn,
    input          i_valid,
    output         o_ready,
    input   [31:0] i_data,
    output  [31:0] o_data
);

endmodule

